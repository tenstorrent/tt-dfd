// SPDX-FileCopyrightText: Copyright 2025 Tenstorrent AI ULC
// SPDX-License-Identifier: Apache-2.0

package mem_gen_pkg;
typedef enum int {
mem_cell_undefined
} MemCell_e;
endpackage : mem_gen_pkg
