package mem_gen_pkg;
typedef enum int {
mem_cell_undefined
} MemCell_e;
endpackage : mem_gen_pkg
