//Include packages below

